interface iface(input logic clk,rst);
   logic WREQ,RREQ;
   logic [7:0] WD,RD;
   logic       e,f;
   
endinterface
